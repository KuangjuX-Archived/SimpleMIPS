module cache(
    input clk_i

);

endmodule: cache